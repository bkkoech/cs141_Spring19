`timescale 1ns / 1ps
`default_nettype none //helps catch typo-related bugs
//////////////////////////////////////////////////////////////////////////////////
// 
// CS 141 - Fall 2015
// Module Name:    and 
// Author(s): 
// Description: 
//
//
//////////////////////////////////////////////////////////////////////////////////
module and(X,Y,Z);

	//parameter definitions
	input wire X[31:0]
	input wire Y[31:0]

	//port definitions - customize for different bit widths


endmodule
`default_nettype wire //some Xilinx IP requires that the default_nettype be set to wire
