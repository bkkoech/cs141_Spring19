`timescale 1ns / 1ps
`default_nettype none //helps catch typo-related bugs
//////////////////////////////////////////////////////////////////////////////////
// 
// CS 141 - Fall 2015
// Module Name:    logical_shifter 
// Author(s): 
// Description: 
//
//
//////////////////////////////////////////////////////////////////////////////////
module logical_shifter();

	//parameter definitions

	//port definitions - customize for different bit widths


endmodule
`default_nettype wire //some Xilinx IP requires that the default_nettype be set to wire
