`timescale 1ns / 1ps
`default_nettype none //helps catch typo-related bugs
//////////////////////////////////////////////////////////////////////////////////
// 
// CS 141 - Fall 2015
// Module Name:    logical_shift_right 
// Author(s): 
// Description: 
//
//
//////////////////////////////////////////////////////////////////////////////////
module logical_shift_right();

// make later
	


endmodule
`default_nettype wire //some Xilinx IP requires that the default_nettype be set to wire
